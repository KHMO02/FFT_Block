class transaction;
logic clk;
logic rst_n; 
logic [11:0] x_r;   
logic [11:0] x_i;   
logic [11:0] X_r;   
logic [11:0] X_i;   
endclass //transaction