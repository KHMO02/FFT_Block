package pack;

`include "transaction.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "sequencer.sv"
`include "subscriber.sv"
`include "env.sv"

    
endpackage